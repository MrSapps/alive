Example VH file :)